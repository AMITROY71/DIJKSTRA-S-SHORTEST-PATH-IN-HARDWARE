`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    19:58:59 01/29/2020 
// Design Name: 
// Module Name:    prom 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module prom_DMH(

input wire [3:0] addr,
input wire [7:0] key_code,
output reg [0:31] M
    );

reg [0:31] rom_A [0:15];
reg [0:31] rom_B [0:15];
reg [0:31] rom_C [0:15];
reg [0:31] rom_D [0:15];
reg [0:31] rom_E [0:15];
reg [0:31] rom_F [0:15];
reg [0:31] rom_G [0:15];
reg [0:31] rom_H [0:15];
reg [0:31] rom_I [0:15];
reg [0:31] rom_J [0:15];
reg [0:31] rom_K [0:15];
reg [0:31] rom_L [0:15];
reg [0:31] rom_M [0:15];
reg [0:31] rom_N [0:15];
reg [0:31] rom_O [0:15];
reg [0:31] rom_P [0:15];
reg [0:31] rom_Q [0:15];
reg [0:31] rom_R [0:15];
reg [0:31] rom_S [0:15];
reg [0:31] rom_T [0:15];
reg [0:31] rom_U [0:15];
reg [0:31] rom_V [0:15];
reg [0:31] rom_W [0:15];
reg [0:31] rom_X [0:15];
reg [0:31] rom_Y [0:15];
reg [0:31] rom_Z [0:15];
reg [0:31] rom_white [0:15];

parameter data_A = {

							32'b00000000000000000000000000000000,
							32'b00000000000000000000000000000000,
							32'b00000000000000000000000000111000,
							32'b00000000000000000000000001101100,
							32'b00000000000000000000000011000110,
							32'b00000000000000000000000011000110,
							32'b00000000000000000000000011000110,
							32'b00000000000000000000000011111110,
							32'b00000000000000000000000011000110,
							32'b00000000000000000000000011000110,
							32'b00000000000000000000000011000110,
							32'b00000000000000000000000011000110,
							32'b00000000000000000000000000000000,
							32'b00000000000000000000000000000000,
							32'b00000000000000000000000000000000,
							32'b00000000000000000000000000000000
	                        
	};                      
	                        
	parameter data_B = {    
                            
							32'b00000000000000000000000000000000,
							32'b00000000000000000000000000000000,
							32'b00000000000000000000000011111100,
							32'b00000000000000000000000001100110,
							32'b00000000000000000000000001100110,
							32'b00000000000000000000000001100110,
							32'b00000000000000000000000001111100,
							32'b00000000000000000000000001100110,
							32'b00000000000000000000000001100110,
							32'b00000000000000000000000001100110,
							32'b00000000000000000000000001100110,
							32'b00000000000000000000000011111100,
							32'b00000000000000000000000000000000,
							32'b00000000000000000000000000000000,
							32'b00000000000000000000000000000000,
							32'b00000000000000000000000000000000
	                        
	};                      
	                        
	parameter data_C = {    
                            
							32'b00000000000000000000000000000000,
							32'b00000000000000000000000000000000,
							32'b00000000000000000000000001111100,
							32'b00000000000000000000000011000110,
							32'b00000000000000000000000011000110,
							32'b00000000000000000000000011000000,
							32'b00000000000000000000000011000000,
							32'b00000000000000000000000011000000,
							32'b00000000000000000000000011000000,
							32'b00000000000000000000000011000110,
							32'b00000000000000000000000011000110,
							32'b00000000000000000000000001111100,
							32'b00000000000000000000000000000000,
							32'b00000000000000000000000000000000,
							32'b00000000000000000000000000000000,
							32'b00000000000000000000000000000000
	                        
	};                      
	                        
	parameter data_D = {    
                            
							32'b00000000000000000000000000000000,
							32'b00000000000000000000000000000000,
							32'b00000000000000000000000011111100,
							32'b00000000000000000000000001100110,
							32'b00000000000000000000000001100110,
							32'b00000000000000000000000001100110,
							32'b00000000000000000000000001100110,
							32'b00000000000000000000000001100110,
							32'b00000000000000000000000001100110,
							32'b00000000000000000000000001100110,
							32'b00000000000000000000000001100110,
							32'b00000000000000000000000011111100,
							32'b00000000000000000000000000000000,
							32'b00000000000000000000000000000000,
							32'b00000000000000000000000000000000,
							32'b00000000000000000000000000000000
	                        
	};                      
	                        
	parameter data_E = {    
                            
							32'b00000000000000000000000000000000,
							32'b00000000000000000000000000000000,
							32'b00000000000000000000000011111110,
							32'b00000000000000000000000001100110,
							32'b00000000000000000000000001100010,
							32'b00000000000000000000000001101000,
							32'b00000000000000000000000001111000,
							32'b00000000000000000000000001111000,
							32'b00000000000000000000000001101000,
							32'b00000000000000000000000001100010,
							32'b00000000000000000000000001100110,
							32'b00000000000000000000000011111110,
							32'b00000000000000000000000000000000,
							32'b00000000000000000000000000000000,
							32'b00000000000000000000000000000000,
							32'b00000000000000000000000000000000
	                        
	};                      
	                        
	parameter data_F = {    
                            
							32'b00000000000000000000000000000000,
							32'b00000000000000000000000000000000,
							32'b00000000000000000000000011111110,
							32'b00000000000000000000000001100110,
							32'b00000000000000000000000001100010,
							32'b00000000000000000000000001101000,
							32'b00000000000000000000000001111000,
							32'b00000000000000000000000001111000,
							32'b00000000000000000000000001101000,
							32'b00000000000000000000000001100000,
							32'b00000000000000000000000001100000,
							32'b00000000000000000000000011110000,
							32'b00000000000000000000000000000000,
							32'b00000000000000000000000000000000,
							32'b00000000000000000000000000000000,
							32'b00000000000000000000000000000000
	                        
	};                      
	                        
	parameter data_G = {    
                            
							32'b00000000000000000000000000000000,
							32'b00000000000000000000000000000000,
							32'b00000000000000000000000001111100,
							32'b00000000000000000000000011000110,
							32'b00000000000000000000000011000110,
							32'b00000000000000000000000011000000,
							32'b00000000000000000000000011000000,
							32'b00000000000000000000000011001110,
							32'b00000000000000000000000011000110,
							32'b00000000000000000000000011000110,
							32'b00000000000000000000000011000110,
							32'b00000000000000000000000001111110,
							32'b00000000000000000000000000000000,
							32'b00000000000000000000000000000000,
							32'b00000000000000000000000000000000,
							32'b00000000000000000000000000000000
	                        
	};                      
	                        
	parameter data_H = {    
                            
							32'b00000000000000000000000000000000,
							32'b00000000000000000000000000000000,
							32'b00000000000000000000000011000110,
							32'b00000000000000000000000011000110,
							32'b00000000000000000000000011000110,
							32'b00000000000000000000000011000110,
							32'b00000000000000000000000011111110,
							32'b00000000000000000000000011000110,
							32'b00000000000000000000000011000110,
							32'b00000000000000000000000011000110,
							32'b00000000000000000000000011000110,
							32'b00000000000000000000000011000110,
							32'b00000000000000000000000000000000,
							32'b00000000000000000000000000000000,
							32'b00000000000000000000000000000000,
							32'b00000000000000000000000000000000
	                        
	};                      
	                        
	parameter data_I = {    
                            
							32'b00000000000000000000000000000000,
							32'b00000000000000000000000000000000,
							32'b00000000000000000000000000111100,
							32'b00000000000000000000000000011000,
							32'b00000000000000000000000000011000,
							32'b00000000000000000000000000011000,
							32'b00000000000000000000000000011000,
							32'b00000000000000000000000000011000,
							32'b00000000000000000000000000011000,
							32'b00000000000000000000000000011000,
							32'b00000000000000000000000000011000,
							32'b00000000000000000000000000111100,
							32'b00000000000000000000000000000000,
							32'b00000000000000000000000000000000,
							32'b00000000000000000000000000000000,
							32'b00000000000000000000000000000000
	                        
	};                      
	                        
	parameter data_J = {    
                            
							32'b00000000000000000000000000000000,
							32'b00000000000000000000000000000000,
							32'b00000000000000000000000000011110,
							32'b00000000000000000000000000001100,
							32'b00000000000000000000000000001100,
							32'b00000000000000000000000000001100,
							32'b00000000000000000000000000001100,
							32'b00000000000000000000000000001100,
							32'b00000000000000000000000011001100,
							32'b00000000000000000000000011001100,
							32'b00000000000000000000000011001100,
							32'b00000000000000000000000001111000,
							32'b00000000000000000000000000000000,
							32'b00000000000000000000000000000000,
							32'b00000000000000000000000000000000,
							32'b00000000000000000000000000000000
	                        
	};                      
	                        
	parameter data_K = {    
                            
							32'b00000000000000000000000000000000,
							32'b00000000000000000000000000000000,
							32'b00000000000000000000000011100110,
							32'b00000000000000000000000001100110,
							32'b00000000000000000000000001100110,
							32'b00000000000000000000000001101100,
							32'b00000000000000000000000001111000,
							32'b00000000000000000000000001111000,
							32'b00000000000000000000000001101100,
							32'b00000000000000000000000001100110,
							32'b00000000000000000000000001100110,
							32'b00000000000000000000000011100110,
							32'b00000000000000000000000000000000,
							32'b00000000000000000000000000000000,
							32'b00000000000000000000000000000000,
							32'b00000000000000000000000000000000
	                        
	};                      
	                        
	parameter data_L = {    
                            
							32'b00000000000000000000000000000000,
							32'b00000000000000000000000000000000,
							32'b00000000000000000000000011110000,
							32'b00000000000000000000000001100000,
							32'b00000000000000000000000001100000,
							32'b00000000000000000000000001100000,
							32'b00000000000000000000000001100000,
							32'b00000000000000000000000001100000,
							32'b00000000000000000000000001100000,
							32'b00000000000000000000000001100010,
							32'b00000000000000000000000001100110,
							32'b00000000000000000000000011111110,
							32'b00000000000000000000000000000000,
							32'b00000000000000000000000000000000,
							32'b00000000000000000000000000000000,
							32'b00000000000000000000000000000000
	                        
	};                      
	                        
	parameter data_M = {    
                            
							32'b00000000000000000000000000000000,
							32'b00000000000000000000000000000000,
							32'b00000000000000000000000010000010,
							32'b00000000000000000000000011000110,
							32'b00000000000000000000000011101110,
							32'b00000000000000000000000011111110,
							32'b00000000000000000000000011111110,
							32'b00000000000000000000000011010110,
							32'b00000000000000000000000011000110,
							32'b00000000000000000000000011000110,
							32'b00000000000000000000000011000110,
							32'b00000000000000000000000011000110,
							32'b00000000000000000000000000000000,
							32'b00000000000000000000000000000000,
							32'b00000000000000000000000000000000,
							32'b00000000000000000000000000000000
	                        
	};                      
	                        
	parameter data_N = {    
                            
							32'b00000000000000000000000000000000,
							32'b00000000000000000000000000000000,
							32'b00000000000000000000000010000110,
							32'b00000000000000000000000011000110,
							32'b00000000000000000000000011100110,
							32'b00000000000000000000000011110110,
							32'b00000000000000000000000011111110,
							32'b00000000000000000000000011011110,
							32'b00000000000000000000000011001110,
							32'b00000000000000000000000011000110,
							32'b00000000000000000000000011000110,
							32'b00000000000000000000000011000110,
							32'b00000000000000000000000000000000,
							32'b00000000000000000000000000000000,
							32'b00000000000000000000000000000000,
							32'b00000000000000000000000000000000
	                        
	};                      
	                        
	parameter data_O = {    
                            
							32'b00000000000000000000000000000000,
							32'b00000000000000000000000000000000,
							32'b00000000000000000000000001111100,
							32'b00000000000000000000000011000110,
							32'b00000000000000000000000011000110,
							32'b00000000000000000000000011000110,
							32'b00000000000000000000000011000110,
							32'b00000000000000000000000011000110,
							32'b00000000000000000000000011000110,
							32'b00000000000000000000000011000110,
							32'b00000000000000000000000011000110,
							32'b00000000000000000000000001111100,
							32'b00000000000000000000000000000000,
							32'b00000000000000000000000000000000,
							32'b00000000000000000000000000000000,
							32'b00000000000000000000000000000000
	                        
	};                      
	                        
	parameter data_P = {    
                            
							32'b00000000000000000000000000000000,
							32'b00000000000000000000000000000000,
							32'b00000000000000000000000011111100,
							32'b00000000000000000000000001100110,
							32'b00000000000000000000000001100110,
							32'b00000000000000000000000001100110,
							32'b00000000000000000000000001100110,
							32'b00000000000000000000000001111100,
							32'b00000000000000000000000001100000,
							32'b00000000000000000000000001100000,
							32'b00000000000000000000000001100000,
							32'b00000000000000000000000011110000,
							32'b00000000000000000000000000000000,
							32'b00000000000000000000000000000000,
							32'b00000000000000000000000000000000,
							32'b00000000000000000000000000000000
	                        
	};                      
	                        
	parameter data_Q = {    
                            
							32'b00000000000000000000000000000000,
							32'b00000000000000000000000000000000,
							32'b00000000000000000000000001111100,
							32'b00000000000000000000000011000110,
							32'b00000000000000000000000011000110,
							32'b00000000000000000000000011000110,
							32'b00000000000000000000000011000110,
							32'b00000000000000000000000011000110,
							32'b00000000000000000000000011000110,
							32'b00000000000000000000000011010110,
							32'b00000000000000000000000011011110,
							32'b00000000000000000000000001111100,
							32'b00000000000000000000000000000110,
							32'b00000000000000000000000000000000,
							32'b00000000000000000000000000000000,
							32'b00000000000000000000000000000000
	                        
	};                      
	                        
	parameter data_R = {    
                            
							32'b00000000000000000000000000000000,
							32'b00000000000000000000000000000000,
							32'b00000000000000000000000011111100,
							32'b00000000000000000000000001100110,
							32'b00000000000000000000000001100110,
							32'b00000000000000000000000001100110,
							32'b00000000000000000000000001100110,
							32'b00000000000000000000000001111100,
							32'b00000000000000000000000001101100,
							32'b00000000000000000000000001100110,
							32'b00000000000000000000000001100110,
							32'b00000000000000000000000011100110,
							32'b00000000000000000000000000000000,
							32'b00000000000000000000000000000000,
							32'b00000000000000000000000000000000,
							32'b00000000000000000000000000000000
	                        
	};                      
	                        
	parameter data_S = {    
                            
							32'b00000000000000000000000000000000,
							32'b00000000000000000000000000000000,
							32'b00000000000000000000000001111100,
							32'b00000000000000000000000011000110,
							32'b00000000000000000000000011000110,
							32'b00000000000000000000000001100000,
							32'b00000000000000000000000000111000,
							32'b00000000000000000000000000001100,
							32'b00000000000000000000000000000110,
							32'b00000000000000000000000011000110,
							32'b00000000000000000000000011000110,
							32'b00000000000000000000000001111100,
							32'b00000000000000000000000000000000,
							32'b00000000000000000000000000000000,
							32'b00000000000000000000000000000000,
							32'b00000000000000000000000000000000
	                        
	};                      
	                        
	parameter data_T = {    
                            
							32'b00000000000000000000000000000000,
							32'b00000000000000000000000000000000,
							32'b00000000000000000000000001111110,
							32'b00000000000000000000000001111110,
							32'b00000000000000000000000001011010,
							32'b00000000000000000000000000011000,
							32'b00000000000000000000000000011000,
							32'b00000000000000000000000000011000,
							32'b00000000000000000000000000011000,
							32'b00000000000000000000000000011000,
							32'b00000000000000000000000000011000,
							32'b00000000000000000000000000111100,
							32'b00000000000000000000000000000000,
							32'b00000000000000000000000000000000,
							32'b00000000000000000000000000000000,
							32'b00000000000000000000000000000000
	                        
	};                      
	                        
	parameter data_U = {    
                            
							32'b00000000000000000000000000000000,
							32'b00000000000000000000000000000000,
							32'b00000000000000000000000011000110,
							32'b00000000000000000000000011000110,
							32'b00000000000000000000000011000110,
							32'b00000000000000000000000011000110,
							32'b00000000000000000000000011000110,
							32'b00000000000000000000000011000110,
							32'b00000000000000000000000011000110,
							32'b00000000000000000000000011000110,
							32'b00000000000000000000000011000110,
							32'b00000000000000000000000001111100,
							32'b00000000000000000000000000000000,
							32'b00000000000000000000000000000000,
							32'b00000000000000000000000000000000,
							32'b00000000000000000000000000000000
	                        
	};                      
	                        
	parameter data_V = {    
                            
							32'b00000000000000000000000000000000,
							32'b00000000000000000000000000000000,
							32'b00000000000000000000000011000110,
							32'b00000000000000000000000011000110,
							32'b00000000000000000000000011000110,
							32'b00000000000000000000000011000110,
							32'b00000000000000000000000011000110,
							32'b00000000000000000000000011000110,
							32'b00000000000000000000000011000110,
							32'b00000000000000000000000001101100,
							32'b00000000000000000000000000111000,
							32'b00000000000000000000000000010000,
							32'b00000000000000000000000000000000,
							32'b00000000000000000000000000000000,
							32'b00000000000000000000000000000000,
							32'b00000000000000000000000000000000
	                        
	};                      
	                        
	parameter data_W = {    
                            
							32'b00000000000000000000000000000000,
							32'b00000000000000000000000000000000,
							32'b00000000000000000000000011000110,
							32'b00000000000000000000000011000110,
							32'b00000000000000000000000011000110,
							32'b00000000000000000000000011000110,
							32'b00000000000000000000000011000110,
							32'b00000000000000000000000011010110,
							32'b00000000000000000000000011111110,
							32'b00000000000000000000000011101110,
							32'b00000000000000000000000011000110,
							32'b00000000000000000000000010000010,
							32'b00000000000000000000000000000000,
							32'b00000000000000000000000000000000,
							32'b00000000000000000000000000000000,
							32'b00000000000000000000000000000000
	                        
	};                      
	                        
	parameter data_X = {    
                            
							32'b00000000000000000000000000000000,
							32'b00000000000000000000000000000000,
							32'b00000000000000000000000011000110,
							32'b00000000000000000000000011000110,
							32'b00000000000000000000000001101100,
							32'b00000000000000000000000001111100,
							32'b00000000000000000000000000111000,
							32'b00000000000000000000000000111000,
							32'b00000000000000000000000001111100,
							32'b00000000000000000000000001101100,
							32'b00000000000000000000000011000110,
							32'b00000000000000000000000011000110,
							32'b00000000000000000000000000000000,
							32'b00000000000000000000000000000000,
							32'b00000000000000000000000000000000,
							32'b00000000000000000000000000000000
	                        
	};                      
	                        
	parameter data_Y = {    
                            
							32'b00000000000000000000000000000000,
							32'b00000000000000000000000000000000,
							32'b00000000000000000000000001100110,
							32'b00000000000000000000000001100110,
							32'b00000000000000000000000001100110,
							32'b00000000000000000000000001100110,
							32'b00000000000000000000000000111100,
							32'b00000000000000000000000000011000,
							32'b00000000000000000000000000011000,
							32'b00000000000000000000000000011000,
							32'b00000000000000000000000000011000,
							32'b00000000000000000000000000111100,
							32'b00000000000000000000000000000000,
							32'b00000000000000000000000000000000,
							32'b00000000000000000000000000000000,
							32'b00000000000000000000000000000000
	                        
	};                      
	                        
	parameter data_Z = {    
                            
							32'b00000000000000000000000000000000,
							32'b00000000000000000000000000000000,
							32'b00000000000000000000000011111110,
							32'b00000000000000000000000011000110,
							32'b00000000000000000000000010000110,
							32'b00000000000000000000000000001100,
							32'b00000000000000000000000000011000,
							32'b00000000000000000000000000110000,
							32'b00000000000000000000000001100000,
							32'b00000000000000000000000011000010,
							32'b00000000000000000000000011000110,
							32'b00000000000000000000000011111110,
							32'b00000000000000000000000000000000,
							32'b00000000000000000000000000000000,
							32'b00000000000000000000000000000000,
							32'b00000000000000000000000000000000
	
	};
	
	parameter data_white = {

	32'b11111111111111111111111111111111,
	32'b11111111111111111111111111111111,
	32'b11111111111111111111111111111111,
	32'b11111111111111111111111111111111,
	32'b11111111111111111111111111111111,
	32'b11111111111111111111111111111111,
	32'b11111111111111111111111111111111,
	32'b11111111111111111111111111111111,
	32'b11111111111111111111111111111111,
	32'b11111111111111111111111111111111,
	32'b11111111111111111111111111111111,
	32'b11111111111111111111111111111111,
	32'b11111111111111111111111111111111,
	32'b11111111111111111111111111111111,
	32'b11111111111111111111111111111111,
	32'b11111111111111111111111111111111
	
	};
	
	
	integer i;
	
	initial
		begin
			for (i = 0; i < 16; i = i + 1)
				begin
					rom_A [i] = data_A[(511-32*i)-:32];
					rom_B [i] = data_B[(511-32*i)-:32];
					rom_C [i] = data_C[(511-32*i)-:32];
					rom_D [i] = data_D[(511-32*i)-:32];
					rom_E [i] = data_E[(511-32*i)-:32];
					rom_F [i] = data_F[(511-32*i)-:32];
					rom_G [i] = data_G[(511-32*i)-:32];
					rom_H [i] = data_H[(511-32*i)-:32];
					rom_I [i] = data_I[(511-32*i)-:32];
					rom_J [i] = data_J[(511-32*i)-:32];
					rom_K [i] = data_K[(511-32*i)-:32];
					rom_L [i] = data_L[(511-32*i)-:32];
					rom_M [i] = data_M[(511-32*i)-:32];
					rom_N [i] = data_N[(511-32*i)-:32];
					rom_O [i] = data_O[(511-32*i)-:32];
					rom_P [i] = data_P[(511-32*i)-:32];
					rom_Q [i] = data_Q[(511-32*i)-:32];
					rom_R [i] = data_R[(511-32*i)-:32];
					rom_S [i] = data_S[(511-32*i)-:32];
					rom_T [i] = data_T[(511-32*i)-:32];
					rom_U [i] = data_U[(511-32*i)-:32];
					rom_V [i] = data_V[(511-32*i)-:32];
					rom_W [i] = data_W[(511-32*i)-:32];
					rom_X [i] = data_X[(511-32*i)-:32];
					rom_Y [i] = data_Y[(511-32*i)-:32];
					rom_Z [i] = data_Z[(511-32*i)-:32];
					rom_white [i] = data_white[(511-32*i)-:32];					
				end
		end
	
	
	always @(key_code or addr)
		begin
			case (key_code)

				8'h1c:  M  =  rom_A[addr];  //  A 
				8'h32:  M  =  rom_B[addr];  //  B 
				8'h21:  M  =  rom_C[addr];  //  C 
				8'h23:  M  =  rom_D[addr];  //  D 
				8'h24:  M  =  rom_E[addr];  //  E 
				8'h2b:  M  =  rom_F[addr];  //  F 
				8'h34:  M  =  rom_G[addr];  //  G 
				8'h33:  M  =  rom_H[addr];  //  H 
				8'h43:  M  =  rom_I[addr];  //  I 
				8'h3b:  M  =  rom_J[addr];  //  J 
				8'h42:  M  =  rom_K[addr];  //  K 
				8'h4b:  M  =  rom_L[addr];  //  L 
				8'h3a:  M  =  rom_M[addr];  //  M 
				8'h31:  M  =  rom_N[addr];  //  N 
				8'h44:  M  =  rom_O[addr];  //  O 
				8'h4d:  M  =  rom_P[addr];  //  P 
				8'h15:  M  =  rom_Q[addr];  //  Q 
				8'h2d:  M  =  rom_R[addr];  //  R 
				8'h1b:  M  =  rom_S[addr];  //  S 
				8'h2c:  M  =  rom_T[addr];  //  T 
				8'h3c:  M  =  rom_U[addr];  //  U 
				8'h2a:  M  =  rom_V[addr];  //  V 
				8'h1d:  M  =  rom_W[addr];  //  W 
				8'h22:  M  =  rom_X[addr];  //  X 
				8'h35:  M  =  rom_Y[addr];  //  Y 
				8'h1a:  M  =  rom_Z[addr];  //  Z 
	
				default:M  =  rom_white[addr];
			endcase
		end
	

endmodule
